
library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity RISCV_ALU is
port(
		--inputs
	    A      : in std_logic_vector(31 downto 0);
	    B      : in std_logic_vector(31 downto 0);
            ALU_ctrl  : in std_logic_vector(3 downto 0);
		--outputs
            result    : out std_logic_vector(31 downto 0);
	--flags
            overflow  : out std_logic;
            negative  : out std_logic;
            zero      : out std_logic;
	    carry     : out std_logic);

end entity;

architecture behave of RISCV_ALU is
	signal temp_result : std_logic_vector(32 downto 0);
	signal V : std_logic;
begin

	process (ALU_ctrl, A, B) is
	variable inputA : signed(32 downto 0);
	variable inputB : signed(32 downto 0);
	variable shiftNum : integer;
	begin
		inputA := signed('0' & A);
		inputB := signed('0' & B);	
		shiftNum := to_integer(unsigned(B));


		case ALU_ctrl is
			when "0000" => --add
				temp_result <= std_logic_vector(signed('0' & A) + signed('0' & B));

			when "0001" | "0111" | "1000" =>  --sub, slt, sltu. Improvement, re-use the sub hardware.
				temp_result <= std_logic_vector(signed('0' & A) + ('0' & (not signed(B) + 1)));

			when "0010" =>  --and (if it turns out that flags are logical, stop setting output will disallow check).
				temp_result(31 downto 0) <= A and B;

			when "0011" =>  --or
				temp_result(31 downto 0) <= A or B;

			when "0100" =>  --xor
				temp_result(31 downto 0) <= A xor B;

			when "0101" =>  --sll --add #B 0's to left of A (I am aware of built-in function, was just curious).
				if shiftNum /= 0 then

				for i in 31 downto shiftNum loop
				inputA(i) := inputA(i-shiftNum);
				end loop;

				for i in shiftNum-1 downto 0 loop
				inputA(i) := '0';
				end loop;

				end if;
			
				temp_result <= std_logic_vector(inputA);

			when "0110" => --srl --add 0 to right

				if shiftNum /= 0 and shiftNum < 32 then
				for i in 0 to 31-shiftNum loop --opposite direction as to not attempt to grab undefined values.
				inputA(i) := inputA(i+shiftNum);
				end loop;

				for i in 32-shiftNum to 31 loop
				inputA(i) := '0';
				end loop;

				elsif shiftNum >= 32 then
				for i in 0 to 31 loop
				inputA(i) := '0';
				end loop;

				end if;

				temp_result <= std_logic_vector(inputA);

			when "1001" =>  --sra:
				if shiftNum /= 0 and shiftNum < 32 then

				for i in 0 to 31-shiftNum loop --opposite direction as to not attempt to grab undefined values.
				inputA(i) := inputA(i+shiftNum);
				end loop;

				for i in 32-shiftNum to 31 loop
				inputA(i) := inputA(31-shiftNum);
				end loop;
				
				elsif shiftNum >= 32 then
				
				for i in 0 to 31 loop
				inputA(i) := inputA(31);
				end loop;				
				
				end if;

				temp_result <= std_logic_vector(inputA);
				
			when others =>
				temp_result <= (others => '0');
		end case;
	end process;

	process (A, B, Temp_Result, ALU_ctrl)
	begin
		if (ALU_ctrl = "0000") then
		V <= (A(31) and B(31) and not(temp_result(31))) or (not(A(31)) and not(B(31)) and temp_result(31));
		
		else
		
		V <= (A(31) and not(B(31)) and not(temp_result(31))) or (not(A(31)) and B(31) and temp_result(31));
		
		end if;
	end process;
	
	with ALU_ctrl select
	result <= (x"0000000" & "000" & (temp_result(31) xor V)) when "0111", --slt
			  (x"0000000" & "000" & not temp_result(32)) when "1000", --sltu
			   temp_result(31 downto 0) when others;
	
	overflow <= V when alu_ctrl = "0000" or alu_ctrl = "0001" else '0';
	
	zero <= '1' when to_integer(signed(temp_result(31 downto 0))) = 0 else '0';
	
	negative <= temp_result(31) when alu_ctrl = "0000" or ALU_ctrl = "0001" else '0';
	
	carry <= temp_result(32) when ALU_ctrl = "0000" or ALU_ctrl = "0001" else '0';

end architecture;
